`timescale 1ns / 1ps

/*
 * Group_ID-61 (15114031_15114032) - Haresh Khanna & Harjot Singh Oberai
 * Date: October 25, 2016
 * adder8bit.v
 *
 */

module mul8bit(
	input wire [7:0] a,
	input wire [7:0] b,
	output wire [15:0] result
    );


endmodule
